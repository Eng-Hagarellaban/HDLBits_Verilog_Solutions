//we want to assign 1 to the output one.
module top_module( output one );

// Insert your code here
    assign one = 1;

endmodule

